<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-60.8454,120.26,324.727,-76.8631</PageViewport>
<gate>
<ID>1</ID>
<type>AA_AND2</type>
<position>120.5,58</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>DE_TO</type>
<position>231.5,-21</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>3</ID>
<type>HA_JUNC_2</type>
<position>-17.5,8</position>
<input>
<ID>N_in0</ID>3 </input>
<input>
<ID>N_in1</ID>73 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>DE_TO</type>
<position>231.5,-26</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>231.5,-28.5</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>395</ID>
<type>AE_OR2</type>
<position>201.5,86.5</position>
<input>
<ID>IN_0</ID>397 </input>
<input>
<ID>IN_1</ID>375 </input>
<output>
<ID>OUT</ID>402 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>DE_TO</type>
<position>231.5,-23.5</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>396</ID>
<type>DA_FROM</type>
<position>181,105.5</position>
<input>
<ID>IN_0</ID>401 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID TOX</lparam></gate>
<gate>
<ID>7</ID>
<type>DA_FROM</type>
<position>105.5,57</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_1</lparam></gate>
<gate>
<ID>8</ID>
<type>HA_JUNC_2</type>
<position>224,-27.5</position>
<input>
<ID>N_in0</ID>118 </input>
<input>
<ID>N_in1</ID>154 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>-42,8</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>HA_JUNC_2</type>
<position>224,-28.5</position>
<input>
<ID>N_in0</ID>120 </input>
<input>
<ID>N_in1</ID>155 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>400</ID>
<type>AE_OR2</type>
<position>213,91</position>
<input>
<ID>IN_0</ID>401 </input>
<input>
<ID>IN_1</ID>402 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>HA_JUNC_2</type>
<position>224,-29.5</position>
<input>
<ID>N_in0</ID>123 </input>
<input>
<ID>N_in1</ID>156 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>HA_JUNC_2</type>
<position>224,-30.5</position>
<input>
<ID>N_in0</ID>128 </input>
<input>
<ID>N_in1</ID>157 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>402</ID>
<type>DE_TO</type>
<position>9,-46.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>13</ID>
<type>DE_TO</type>
<position>139.5,58</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2R1</lparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>9,18.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK0</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_AND2</type>
<position>-30.5,-8.5</position>
<input>
<ID>IN_0</ID>407 </input>
<input>
<ID>IN_1</ID>406 </input>
<output>
<ID>OUT</ID>325 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-27.5</position>
<input>
<ID>N_in0</ID>168 </input>
<input>
<ID>N_in1</ID>118 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>-38,-7.5</position>
<input>
<ID>IN_0</ID>407 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>16</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-28.5</position>
<input>
<ID>N_in0</ID>167 </input>
<input>
<ID>N_in1</ID>120 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-29.5</position>
<input>
<ID>N_in0</ID>166 </input>
<input>
<ID>N_in1</ID>123 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-30.5</position>
<input>
<ID>N_in0</ID>165 </input>
<input>
<ID>N_in1</ID>128 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>408</ID>
<type>DE_TO</type>
<position>36,-104.5</position>
<input>
<ID>IN_0</ID>413 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_AND2</type>
<position>120.5,51</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>DE_TO</type>
<position>36,-109.5</position>
<input>
<ID>IN_0</ID>414 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RD</lparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>105.5,50</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_2</lparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>139.5,51</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2R2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_RAM_4x4</type>
<position>23,-101</position>
<input>
<ID>ADDRESS_0</ID>37 </input>
<input>
<ID>ADDRESS_1</ID>61 </input>
<input>
<ID>ADDRESS_2</ID>62 </input>
<input>
<ID>ADDRESS_3</ID>63 </input>
<input>
<ID>DATA_IN_0</ID>174 </input>
<input>
<ID>DATA_IN_1</ID>175 </input>
<input>
<ID>DATA_IN_2</ID>176 </input>
<input>
<ID>DATA_IN_3</ID>177 </input>
<output>
<ID>DATA_OUT_0</ID>174 </output>
<output>
<ID>DATA_OUT_1</ID>175 </output>
<output>
<ID>DATA_OUT_2</ID>176 </output>
<output>
<ID>DATA_OUT_3</ID>177 </output>
<input>
<ID>ENABLE_0</ID>414 </input>
<input>
<ID>write_clock</ID>152 </input>
<input>
<ID>write_enable</ID>413 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:1 2</lparam>
<lparam>Address:2 3</lparam>
<lparam>Address:3 9</lparam>
<lparam>Address:4 9</lparam>
<lparam>Address:5 2</lparam>
<lparam>Address:6 11</lparam>
<lparam>Address:7 1</lparam>
<lparam>Address:8 1</lparam>
<lparam>Address:9 2</lparam>
<lparam>Address:10 3</lparam>
<lparam>Address:11 5</lparam>
<lparam>Address:12 8</lparam>
<lparam>Address:13 13</lparam>
<lparam>Address:14 5</lparam>
<lparam>Address:15 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_REGISTER4</type>
<position>-12,13.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<output>
<ID>OUT_1</ID>89 </output>
<output>
<ID>OUT_2</ID>90 </output>
<input>
<ID>clear</ID>104 </input>
<input>
<ID>clock</ID>73 </input>
<input>
<ID>count_enable</ID>116 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>24</ID>
<type>BE_ROM_8x8</type>
<position>54.5,6</position>
<input>
<ID>ADDRESS_0</ID>49 </input>
<input>
<ID>ADDRESS_1</ID>48 </input>
<input>
<ID>ADDRESS_2</ID>47 </input>
<input>
<ID>ADDRESS_3</ID>46 </input>
<input>
<ID>ADDRESS_4</ID>45 </input>
<input>
<ID>ADDRESS_5</ID>44 </input>
<input>
<ID>ADDRESS_6</ID>43 </input>
<input>
<ID>ADDRESS_7</ID>42 </input>
<output>
<ID>DATA_OUT_0</ID>38 </output>
<output>
<ID>DATA_OUT_1</ID>39 </output>
<output>
<ID>DATA_OUT_2</ID>40 </output>
<output>
<ID>DATA_OUT_3</ID>41 </output>
<output>
<ID>DATA_OUT_4</ID>34 </output>
<output>
<ID>DATA_OUT_5</ID>35 </output>
<output>
<ID>DATA_OUT_6</ID>36 </output>
<output>
<ID>DATA_OUT_7</ID>271 </output>
<input>
<ID>ENABLE_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 112</lparam>
<lparam>Address:1 96</lparam>
<lparam>Address:2 80</lparam>
<lparam>Address:3 64</lparam>
<lparam>Address:4 48</lparam>
<lparam>Address:5 32</lparam>
<lparam>Address:6 16</lparam>
<lparam>Address:8 255</lparam>
<lparam>Address:13 130</lparam>
<lparam>Address:127 131</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND2</type>
<position>120.5,44.5</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_REGISTER4</type>
<position>-8,-59</position>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>175 </input>
<input>
<ID>IN_2</ID>176 </input>
<input>
<ID>IN_3</ID>177 </input>
<output>
<ID>OUT_0</ID>9 </output>
<output>
<ID>OUT_1</ID>10 </output>
<output>
<ID>OUT_2</ID>11 </output>
<output>
<ID>OUT_3</ID>12 </output>
<input>
<ID>clock</ID>187 </input>
<input>
<ID>load</ID>20 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>231.5,108</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2A</lparam></gate>
<gate>
<ID>28</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>-1,-63.5</position>
<input>
<ID>ENABLE_0</ID>14 </input>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>12 </input>
<output>
<ID>OUT_0</ID>174 </output>
<output>
<ID>OUT_1</ID>175 </output>
<output>
<ID>OUT_2</ID>176 </output>
<output>
<ID>OUT_3</ID>177 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>29</ID>
<type>DE_TO</type>
<position>9,15.5</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK1</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>2.5,-55</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2D</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>-0.5,-91</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2M</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>-9,-49</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2X</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>105.5,43.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_3</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_OR2</type>
<position>223.5,90</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>DE_TO</type>
<position>231.5,-31.5</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>231.5,-36.5</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>231.5,-39</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>231.5,-34</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>39</ID>
<type>HA_JUNC_2</type>
<position>224,-33.5</position>
<input>
<ID>N_in0</ID>25 </input>
<input>
<ID>N_in1</ID>158 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>HA_JUNC_2</type>
<position>224,-34.5</position>
<input>
<ID>N_in0</ID>26 </input>
<input>
<ID>N_in1</ID>159 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>HA_JUNC_2</type>
<position>224,-35.5</position>
<input>
<ID>N_in0</ID>27 </input>
<input>
<ID>N_in1</ID>160 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>HA_JUNC_2</type>
<position>224,-36.5</position>
<input>
<ID>N_in0</ID>28 </input>
<input>
<ID>N_in1</ID>161 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-33.5</position>
<input>
<ID>N_in0</ID>172 </input>
<input>
<ID>N_in1</ID>25 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-34.5</position>
<input>
<ID>N_in0</ID>171 </input>
<input>
<ID>N_in1</ID>26 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-35.5</position>
<input>
<ID>N_in0</ID>170 </input>
<input>
<ID>N_in1</ID>27 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-36.5</position>
<input>
<ID>N_in0</ID>169 </input>
<input>
<ID>N_in1</ID>28 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>6,-63.5</position>
<input>
<ID>ENABLE_0</ID>33 </input>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>12 </input>
<output>
<ID>OUT_0</ID>178 </output>
<output>
<ID>OUT_1</ID>179 </output>
<output>
<ID>OUT_2</ID>180 </output>
<output>
<ID>OUT_3</ID>182 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>10,-60</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID X2A</lparam></gate>
<gate>
<ID>49</ID>
<type>BE_DECODER_3x8</type>
<position>-4,16</position>
<input>
<ID>ENABLE</ID>116 </input>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>90 </input>
<output>
<ID>OUT_0</ID>103 </output>
<output>
<ID>OUT_1</ID>305 </output>
<output>
<ID>OUT_2</ID>304 </output>
<output>
<ID>OUT_3</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_REGISTER4</type>
<position>65.5,-4.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>36 </input>
<input>
<ID>IN_3</ID>271 </input>
<output>
<ID>OUT_0</ID>60 </output>
<output>
<ID>OUT_1</ID>59 </output>
<output>
<ID>OUT_2</ID>58 </output>
<output>
<ID>OUT_3</ID>57 </output>
<input>
<ID>clear</ID>112 </input>
<input>
<ID>clock</ID>100 </input>
<input>
<ID>load</ID>50 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>139.5,44.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2R3</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_REGISTER4</type>
<position>65.5,-17.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>41 </input>
<output>
<ID>OUT_0</ID>51 </output>
<output>
<ID>OUT_1</ID>52 </output>
<output>
<ID>OUT_2</ID>53 </output>
<output>
<ID>OUT_3</ID>54 </output>
<input>
<ID>clear</ID>112 </input>
<input>
<ID>clock</ID>100 </input>
<input>
<ID>load</ID>50 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_TOGGLE</type>
<position>-28,3.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_REGISTER8</type>
<position>43,5.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>41 </input>
<input>
<ID>IN_4</ID>34 </input>
<input>
<ID>IN_5</ID>35 </input>
<input>
<ID>IN_6</ID>36 </input>
<output>
<ID>OUT_0</ID>49 </output>
<output>
<ID>OUT_1</ID>48 </output>
<output>
<ID>OUT_2</ID>47 </output>
<output>
<ID>OUT_3</ID>46 </output>
<output>
<ID>OUT_4</ID>45 </output>
<output>
<ID>OUT_5</ID>44 </output>
<output>
<ID>OUT_6</ID>43 </output>
<output>
<ID>OUT_7</ID>42 </output>
<input>
<ID>clear</ID>112 </input>
<input>
<ID>clock</ID>318 </input>
<input>
<ID>count_enable</ID>292 </input>
<input>
<ID>load</ID>310 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND2</type>
<position>119.5,98.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>FF_GND</type>
<position>226.5,104.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>72.5,-22</position>
<input>
<ID>ENABLE_0</ID>55 </input>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<input>
<ID>IN_3</ID>54 </input>
<output>
<ID>OUT_0</ID>118 </output>
<output>
<ID>OUT_1</ID>120 </output>
<output>
<ID>OUT_2</ID>123 </output>
<output>
<ID>OUT_3</ID>128 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>76.5,-12.5</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID P2D</lparam></gate>
<gate>
<ID>59</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>79.5,-22</position>
<input>
<ID>ENABLE_0</ID>56 </input>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<input>
<ID>IN_3</ID>54 </input>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>26 </output>
<output>
<ID>OUT_2</ID>27 </output>
<output>
<ID>OUT_3</ID>28 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>84.5,-12.5</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID P2A</lparam></gate>
<gate>
<ID>61</ID>
<type>DE_TO</type>
<position>9.5,3.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RST</lparam></gate>
<gate>
<ID>62</ID>
<type>BI_DECODER_4x16</type>
<position>104,2</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>57 </input>
<output>
<ID>OUT_0</ID>77 </output>
<output>
<ID>OUT_1</ID>78 </output>
<output>
<ID>OUT_2</ID>79 </output>
<output>
<ID>OUT_3</ID>80 </output>
<output>
<ID>OUT_4</ID>81 </output>
<output>
<ID>OUT_5</ID>82 </output>
<output>
<ID>OUT_6</ID>307 </output>
<output>
<ID>OUT_7</ID>308 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>104.5,97.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_REGISTER4</type>
<position>0.5,-101.5</position>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>175 </input>
<input>
<ID>IN_2</ID>176 </input>
<input>
<ID>IN_3</ID>177 </input>
<output>
<ID>OUT_0</ID>67 </output>
<output>
<ID>OUT_1</ID>66 </output>
<output>
<ID>OUT_2</ID>65 </output>
<output>
<ID>OUT_3</ID>64 </output>
<input>
<ID>clock</ID>152 </input>
<input>
<ID>load</ID>24 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_OR2</type>
<position>30.5,-22</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>14.5,-26</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RST</lparam></gate>
<gate>
<ID>67</ID>
<type>BE_DECODER_3x8</type>
<position>154.5,-15</position>
<input>
<ID>ENABLE</ID>153 </input>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<output>
<ID>OUT_0</ID>124 </output>
<output>
<ID>OUT_1</ID>125 </output>
<output>
<ID>OUT_2</ID>126 </output>
<output>
<ID>OUT_3</ID>127 </output>
<output>
<ID>OUT_6</ID>98 </output>
<output>
<ID>OUT_7</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>68</ID>
<type>DA_FROM</type>
<position>167,106</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID MOVEAX</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_OR2</type>
<position>195,76</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>DE_TO</type>
<position>231.5,95</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID P2D</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>173.5,105.5</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID LOADX</lparam></gate>
<gate>
<ID>72</ID>
<type>DE_TO</type>
<position>231.5,99</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2D</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>170,105.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID MOVEXA</lparam></gate>
<gate>
<ID>74</ID>
<type>DE_TO</type>
<position>231.5,76</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID P2A</lparam></gate>
<gate>
<ID>75</ID>
<type>DE_TO</type>
<position>231.5,83.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR</lparam></gate>
<gate>
<ID>76</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>14.5,-94.5</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>179 </input>
<input>
<ID>IN_2</ID>180 </input>
<input>
<ID>IN_3</ID>182 </input>
<output>
<ID>OUT_0</ID>37 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>62 </output>
<output>
<ID>OUT_3</ID>63 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>77</ID>
<type>DE_TO</type>
<position>126.5,20</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID NOP</lparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>124,20</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID LOADX</lparam></gate>
<gate>
<ID>79</ID>
<type>DE_TO</type>
<position>121.5,20</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID XTO</lparam></gate>
<gate>
<ID>80</ID>
<type>DE_TO</type>
<position>119,20</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID TOX</lparam></gate>
<gate>
<ID>81</ID>
<type>DE_TO</type>
<position>116.5,20</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID MOVEXA</lparam></gate>
<gate>
<ID>82</ID>
<type>DE_TO</type>
<position>114,20</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID MOVEAX</lparam></gate>
<gate>
<ID>83</ID>
<type>DE_TO</type>
<position>110,20.5</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID OPER</lparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>112,20</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID IF</lparam></gate>
<gate>
<ID>86</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>7.5,-101</position>
<input>
<ID>ENABLE_0</ID>75 </input>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>66 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>64 </input>
<output>
<ID>OUT_0</ID>37 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>62 </output>
<output>
<ID>OUT_3</ID>63 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>87</ID>
<type>DE_TO</type>
<position>138.5,98.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R12D</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_AND2</type>
<position>119.5,85.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>104.5,84.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_3</lparam></gate>
<gate>
<ID>90</ID>
<type>DE_TO</type>
<position>138.5,85.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R32D</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>119.5,91.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>DA_FROM</type>
<position>104.5,90.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_2</lparam></gate>
<gate>
<ID>94</ID>
<type>DE_TO</type>
<position>138.5,91.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R22D</lparam></gate>
<gate>
<ID>95</ID>
<type>DE_TO</type>
<position>9,10</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK_EXE</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>69,3</position>
<gparam>LABEL_TEXT R_I</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AE_OR2</type>
<position>-6,6.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND2</type>
<position>21,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>22,-19.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK1</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_AND4</type>
<position>94,-23</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<input>
<ID>IN_3</ID>54 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>101</ID>
<type>DE_TO</type>
<position>-10,0</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>14.5,-23</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>101,-23</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AD_IS_F</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>4,-94</position>
<gparam>LABEL_TEXT R_M</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>DA_FROM</type>
<position>26,-90</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AD_IS_F</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>70,-10</position>
<gparam>LABEL_TEXT R_P</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AE_SMALL_INVERTER</type>
<position>20.5,-94.5</position>
<input>
<ID>IN_0</ID>75 </input>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>15,-73.5</position>
<gparam>LABEL_TEXT DATA BUS</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>DA_FROM</type>
<position>40.5,-22.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RST</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>14.5,-79.5</position>
<gparam>LABEL_TEXT ADDRESS BUS</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>DA_FROM</type>
<position>149.5,107</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID GOTO</lparam></gate>
<gate>
<ID>113</ID>
<type>DE_TO</type>
<position>95,17.5</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID GOTO</lparam></gate>
<gate>
<ID>119</ID>
<type>DE_TO</type>
<position>229,-43.5</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WR</lparam></gate>
<gate>
<ID>120</ID>
<type>DE_TO</type>
<position>229,-47</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RD</lparam></gate>
<gate>
<ID>121</ID>
<type>DE_TO</type>
<position>172,-18.5</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R_2</lparam></gate>
<gate>
<ID>122</ID>
<type>DE_TO</type>
<position>172,-15.5</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R_3</lparam></gate>
<gate>
<ID>123</ID>
<type>DE_TO</type>
<position>172,-23.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R_0</lparam></gate>
<gate>
<ID>124</ID>
<type>DE_TO</type>
<position>172,-21</position>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R_1</lparam></gate>
<gate>
<ID>125</ID>
<type>DE_TO</type>
<position>172.5,-8</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R_M</lparam></gate>
<gate>
<ID>126</ID>
<type>DE_TO</type>
<position>172.5,-5.5</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R_Y</lparam></gate>
<gate>
<ID>127</ID>
<type>EE_VDD</type>
<position>-12,22.5</position>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_LABEL</type>
<position>-5,-51</position>
<gparam>LABEL_TEXT R_X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_REGISTER4</type>
<position>69,-59</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>136 </input>
<input>
<ID>IN_2</ID>137 </input>
<input>
<ID>IN_3</ID>138 </input>
<output>
<ID>OUT_0</ID>130 </output>
<output>
<ID>OUT_1</ID>131 </output>
<output>
<ID>OUT_2</ID>132 </output>
<output>
<ID>OUT_3</ID>133 </output>
<input>
<ID>clock</ID>187 </input>
<input>
<ID>load</ID>141 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>131</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>76,-63.5</position>
<input>
<ID>ENABLE_0</ID>134 </input>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>131 </input>
<input>
<ID>IN_2</ID>132 </input>
<input>
<ID>IN_3</ID>133 </input>
<output>
<ID>OUT_0</ID>174 </output>
<output>
<ID>OUT_1</ID>175 </output>
<output>
<ID>OUT_2</ID>176 </output>
<output>
<ID>OUT_3</ID>177 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>79.5,-55</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Y2D</lparam></gate>
<gate>
<ID>133</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>62,-64.5</position>
<input>
<ID>ENABLE_0</ID>139 </input>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>175 </input>
<input>
<ID>IN_2</ID>176 </input>
<input>
<ID>IN_3</ID>177 </input>
<output>
<ID>OUT_0</ID>135 </output>
<output>
<ID>OUT_1</ID>136 </output>
<output>
<ID>OUT_2</ID>137 </output>
<output>
<ID>OUT_3</ID>138 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>58,-60</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2Y</lparam></gate>
<gate>
<ID>135</ID>
<type>HA_JUNC_2</type>
<position>-21,-74.5</position>
<input>
<ID>N_in0</ID>168 </input>
<input>
<ID>N_in1</ID>174 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>HA_JUNC_2</type>
<position>-21,-75.5</position>
<input>
<ID>N_in0</ID>167 </input>
<input>
<ID>N_in1</ID>175 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>64,-52.5</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_Y</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>70,-50.5</position>
<gparam>LABEL_TEXT R_Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>HA_JUNC_2</type>
<position>-21,-76.5</position>
<input>
<ID>N_in0</ID>166 </input>
<input>
<ID>N_in1</ID>176 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AE_FULLADDER_4BIT</type>
<position>23,-60</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>12 </input>
<input>
<ID>IN_B_0</ID>130 </input>
<input>
<ID>IN_B_1</ID>131 </input>
<input>
<ID>IN_B_2</ID>132 </input>
<input>
<ID>IN_B_3</ID>133 </input>
<output>
<ID>OUT_0</ID>145 </output>
<output>
<ID>OUT_1</ID>144 </output>
<output>
<ID>OUT_2</ID>143 </output>
<output>
<ID>OUT_3</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>141</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>23,-67.5</position>
<input>
<ID>ENABLE_0</ID>146 </input>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_2</ID>144 </input>
<input>
<ID>IN_3</ID>145 </input>
<output>
<ID>OUT_0</ID>177 </output>
<output>
<ID>OUT_1</ID>176 </output>
<output>
<ID>OUT_2</ID>175 </output>
<output>
<ID>OUT_3</ID>174 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>32.5,-63.5</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID AD2D</lparam></gate>
<gate>
<ID>144</ID>
<type>HA_JUNC_2</type>
<position>224,-40</position>
<input>
<ID>N_in0</ID>151 </input>
<input>
<ID>N_in1</ID>162 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>HA_JUNC_2</type>
<position>224,-41</position>
<input>
<ID>N_in0</ID>150 </input>
<input>
<ID>N_in1</ID>163 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-40</position>
<input>
<ID>N_in1</ID>151 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>HA_JUNC_2</type>
<position>-18.5,-41</position>
<input>
<ID>N_in1</ID>150 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>HA_JUNC_2</type>
<position>-21,-77.5</position>
<input>
<ID>N_in0</ID>165 </input>
<input>
<ID>N_in1</ID>177 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>DA_FROM</type>
<position>45.5,-99.5</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID CLK_EXE</lparam></gate>
<gate>
<ID>150</ID>
<type>DE_TO</type>
<position>231.5,72.5</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RD</lparam></gate>
<gate>
<ID>151</ID>
<type>HA_JUNC_2</type>
<position>-21,-80.5</position>
<input>
<ID>N_in0</ID>172 </input>
<input>
<ID>N_in1</ID>178 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AE_OR2</type>
<position>147,-11.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>HA_JUNC_2</type>
<position>-21,-81.5</position>
<input>
<ID>N_in0</ID>171 </input>
<input>
<ID>N_in1</ID>179 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>HA_JUNC_2</type>
<position>-21,-82.5</position>
<input>
<ID>N_in0</ID>170 </input>
<input>
<ID>N_in1</ID>180 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>HA_JUNC_2</type>
<position>-21,-83.5</position>
<input>
<ID>N_in0</ID>169 </input>
<input>
<ID>N_in1</ID>182 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>HA_JUNC_2</type>
<position>81.5,-74.5</position>
<input>
<ID>N_in0</ID>174 </input>
<input>
<ID>N_in1</ID>209 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>HA_JUNC_2</type>
<position>81.5,-75.5</position>
<input>
<ID>N_in0</ID>175 </input>
<input>
<ID>N_in1</ID>210 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>HA_JUNC_2</type>
<position>81.5,-76.5</position>
<input>
<ID>N_in0</ID>176 </input>
<input>
<ID>N_in1</ID>211 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>HA_JUNC_2</type>
<position>81.5,-77.5</position>
<input>
<ID>N_in0</ID>177 </input>
<input>
<ID>N_in1</ID>212 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>43,-26</position>
<gparam>LABEL_TEXT DATA BUS</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>42.5,-32</position>
<gparam>LABEL_TEXT ADDRESS BUS</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>118.5,-73.5</position>
<gparam>LABEL_TEXT DATA BUS</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>118,-79.5</position>
<gparam>LABEL_TEXT ADDRESS BUS</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>HA_JUNC_2</type>
<position>81.5,-80.5</position>
<input>
<ID>N_in0</ID>178 </input>
<input>
<ID>N_in1</ID>140 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>HA_JUNC_2</type>
<position>81.5,-81.5</position>
<input>
<ID>N_in0</ID>179 </input>
<input>
<ID>N_in1</ID>148 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>HA_JUNC_2</type>
<position>81.5,-82.5</position>
<input>
<ID>N_in0</ID>180 </input>
<input>
<ID>N_in1</ID>149 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>HA_JUNC_2</type>
<position>81.5,-83.5</position>
<input>
<ID>N_in0</ID>182 </input>
<input>
<ID>N_in1</ID>164 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>DE_TO</type>
<position>232,62</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AD2D</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>161.5,106</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>175</ID>
<type>DE_TO</type>
<position>138,112</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2D</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>103.5,115</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID TOX</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND2</type>
<position>119.5,112</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>186 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>DA_FROM</type>
<position>104,110</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_Y</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_REGISTER4</type>
<position>187,-59</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>210 </input>
<input>
<ID>IN_2</ID>211 </input>
<input>
<ID>IN_3</ID>212 </input>
<output>
<ID>OUT_0</ID>188 </output>
<output>
<ID>OUT_1</ID>189 </output>
<output>
<ID>OUT_2</ID>190 </output>
<output>
<ID>OUT_3</ID>191 </output>
<input>
<ID>clock</ID>187 </input>
<input>
<ID>load</ID>198 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 13</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>182</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>194,-63.5</position>
<input>
<ID>ENABLE_0</ID>192 </input>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>189 </input>
<input>
<ID>IN_2</ID>190 </input>
<input>
<ID>IN_3</ID>191 </input>
<output>
<ID>OUT_0</ID>209 </output>
<output>
<ID>OUT_1</ID>210 </output>
<output>
<ID>OUT_2</ID>211 </output>
<output>
<ID>OUT_3</ID>212 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>183</ID>
<type>DA_FROM</type>
<position>197.5,-55</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID R32D</lparam></gate>
<gate>
<ID>185</ID>
<type>DA_FROM</type>
<position>181.5,-49.5</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2R3</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>188,-50.5</position>
<gparam>LABEL_TEXT R_3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>EE_VDD</type>
<position>60.5,16.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>192</ID>
<type>HA_JUNC_2</type>
<position>206,-74.5</position>
<input>
<ID>N_in0</ID>209 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>193</ID>
<type>HA_JUNC_2</type>
<position>206,-75.5</position>
<input>
<ID>N_in0</ID>210 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>HA_JUNC_2</type>
<position>206,-76.5</position>
<input>
<ID>N_in0</ID>211 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>HA_JUNC_2</type>
<position>206,-77.5</position>
<input>
<ID>N_in0</ID>212 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>HA_JUNC_2</type>
<position>206,-80.5</position>
<input>
<ID>N_in0</ID>140 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>HA_JUNC_2</type>
<position>206,-81.5</position>
<input>
<ID>N_in0</ID>148 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>HA_JUNC_2</type>
<position>206,-82.5</position>
<input>
<ID>N_in0</ID>149 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>HA_JUNC_2</type>
<position>206,-83.5</position>
<input>
<ID>N_in0</ID>164 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>DA_FROM</type>
<position>201,-72</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID CLK_EXE</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_REGISTER4</type>
<position>158.5,-58.5</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>210 </input>
<input>
<ID>IN_2</ID>211 </input>
<input>
<ID>IN_3</ID>212 </input>
<output>
<ID>OUT_0</ID>214 </output>
<output>
<ID>OUT_1</ID>215 </output>
<output>
<ID>OUT_2</ID>216 </output>
<output>
<ID>OUT_3</ID>217 </output>
<input>
<ID>clock</ID>187 </input>
<input>
<ID>load</ID>224 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>210</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>165.5,-63</position>
<input>
<ID>ENABLE_0</ID>218 </input>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>215 </input>
<input>
<ID>IN_2</ID>216 </input>
<input>
<ID>IN_3</ID>217 </input>
<output>
<ID>OUT_0</ID>209 </output>
<output>
<ID>OUT_1</ID>210 </output>
<output>
<ID>OUT_2</ID>211 </output>
<output>
<ID>OUT_3</ID>212 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>211</ID>
<type>DA_FROM</type>
<position>169,-54.5</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID R22D</lparam></gate>
<gate>
<ID>213</ID>
<type>DA_FROM</type>
<position>153,-49.5</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2R2</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>159.5,-50</position>
<gparam>LABEL_TEXT R_2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>AA_REGISTER4</type>
<position>131.5,-58</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>210 </input>
<input>
<ID>IN_2</ID>211 </input>
<input>
<ID>IN_3</ID>212 </input>
<output>
<ID>OUT_0</ID>229 </output>
<output>
<ID>OUT_1</ID>230 </output>
<output>
<ID>OUT_2</ID>231 </output>
<output>
<ID>OUT_3</ID>232 </output>
<input>
<ID>clock</ID>187 </input>
<input>
<ID>load</ID>239 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 11</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>217</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>138.5,-62.5</position>
<input>
<ID>ENABLE_0</ID>233 </input>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>230 </input>
<input>
<ID>IN_2</ID>231 </input>
<input>
<ID>IN_3</ID>232 </input>
<output>
<ID>OUT_0</ID>209 </output>
<output>
<ID>OUT_1</ID>210 </output>
<output>
<ID>OUT_2</ID>211 </output>
<output>
<ID>OUT_3</ID>212 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>142,-54</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID R12D</lparam></gate>
<gate>
<ID>220</ID>
<type>DA_FROM</type>
<position>130.5,-49</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2R1</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>135,-50</position>
<gparam>LABEL_TEXT R_1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_REGISTER4</type>
<position>104.5,-58</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>210 </input>
<input>
<ID>IN_2</ID>211 </input>
<input>
<ID>IN_3</ID>212 </input>
<output>
<ID>OUT_0</ID>244 </output>
<output>
<ID>OUT_1</ID>245 </output>
<output>
<ID>OUT_2</ID>246 </output>
<output>
<ID>OUT_3</ID>247 </output>
<input>
<ID>clock</ID>187 </input>
<input>
<ID>load</ID>254 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 10</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>224</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>111.5,-62.5</position>
<input>
<ID>ENABLE_0</ID>248 </input>
<input>
<ID>IN_0</ID>244 </input>
<input>
<ID>IN_1</ID>245 </input>
<input>
<ID>IN_2</ID>246 </input>
<input>
<ID>IN_3</ID>247 </input>
<output>
<ID>OUT_0</ID>209 </output>
<output>
<ID>OUT_1</ID>210 </output>
<output>
<ID>OUT_2</ID>211 </output>
<output>
<ID>OUT_3</ID>212 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>225</ID>
<type>DA_FROM</type>
<position>115,-54</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID R02D</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>103.5,-49</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2R0</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_LABEL</type>
<position>107.5,-50</position>
<gparam>LABEL_TEXT R_0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>230</ID>
<type>AA_AND2</type>
<position>120.5,37</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>226 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>231</ID>
<type>DA_FROM</type>
<position>105.5,36</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_M</lparam></gate>
<gate>
<ID>232</ID>
<type>DE_TO</type>
<position>139.5,37</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2M</lparam></gate>
<gate>
<ID>247</ID>
<type>AA_AND2</type>
<position>119.5,104.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>259 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>104.5,103.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_0</lparam></gate>
<gate>
<ID>250</ID>
<type>DE_TO</type>
<position>138.5,104.5</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R02D</lparam></gate>
<gate>
<ID>252</ID>
<type>DE_TO</type>
<position>139,74</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2Y</lparam></gate>
<gate>
<ID>253</ID>
<type>DA_FROM</type>
<position>104.5,77</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID XTO</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_AND2</type>
<position>120.5,74</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>263 </input>
<output>
<ID>OUT</ID>261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>DA_FROM</type>
<position>105,72</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_Y</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_AND2</type>
<position>120.5,66.5</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>264 </input>
<output>
<ID>OUT</ID>265 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>DA_FROM</type>
<position>105.5,65.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID R_0</lparam></gate>
<gate>
<ID>258</ID>
<type>DE_TO</type>
<position>139.5,66.5</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2R0</lparam></gate>
<gate>
<ID>259</ID>
<type>DA_FROM</type>
<position>177.5,105.5</position>
<input>
<ID>IN_0</ID>368 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID XTO</lparam></gate>
<gate>
<ID>260</ID>
<type>DA_FROM</type>
<position>42,21.5</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC</lparam></gate>
<gate>
<ID>261</ID>
<type>AE_OR2</type>
<position>191,99</position>
<input>
<ID>IN_0</ID>368 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>262</ID>
<type>DE_TO</type>
<position>231.5,90</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2X</lparam></gate>
<gate>
<ID>265</ID>
<type>DE_TO</type>
<position>232,36</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC</lparam></gate>
<gate>
<ID>289</ID>
<type>EE_VDD</type>
<position>43,19</position>
<output>
<ID>OUT_0</ID>292 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>300</ID>
<type>BB_CLOCK</type>
<position>-27.5,8</position>
<output>
<ID>CLK</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>301</ID>
<type>DE_TO</type>
<position>9,12.5</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK_EXE2</lparam></gate>
<gate>
<ID>304</ID>
<type>DA_FROM</type>
<position>13.5,-11</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK0</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_MUX_2x1</type>
<position>21.5,-9.5</position>
<input>
<ID>IN_0</ID>311 </input>
<input>
<ID>IN_1</ID>313 </input>
<output>
<ID>OUT</ID>314 </output>
<input>
<ID>SEL_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>DA_FROM</type>
<position>18,-5</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RST</lparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>13.5,-8.5</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_OR2</type>
<position>30.5,-11</position>
<input>
<ID>IN_0</ID>314 </input>
<input>
<ID>IN_1</ID>315 </input>
<output>
<ID>OUT</ID>318 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_AND2</type>
<position>22.5,-16</position>
<input>
<ID>IN_0</ID>316 </input>
<input>
<ID>IN_1</ID>317 </input>
<output>
<ID>OUT</ID>315 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>310</ID>
<type>DA_FROM</type>
<position>10.5,-17.5</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK_EXE2</lparam></gate>
<gate>
<ID>311</ID>
<type>DA_FROM</type>
<position>13,-14</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IS_IF</lparam></gate>
<gate>
<ID>313</ID>
<type>DA_FROM</type>
<position>-38,-11</position>
<input>
<ID>IN_0</ID>406 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID IF</lparam></gate>
<gate>
<ID>314</ID>
<type>DA_FROM</type>
<position>-35.5,-14</position>
<input>
<ID>IN_0</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>315</ID>
<type>DE_TO</type>
<position>-9.5,-8.5</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID IS_IF</lparam></gate>
<gate>
<ID>317</ID>
<type>BE_JKFF_LOW</type>
<position>-16.5,-10.5</position>
<input>
<ID>J</ID>325 </input>
<input>
<ID>K</ID>322 </input>
<output>
<ID>Q</ID>319 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>318</ID>
<type>AE_SMALL_INVERTER</type>
<position>-23.5,-12.5</position>
<input>
<ID>IN_0</ID>325 </input>
<output>
<ID>OUT_0</ID>322 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>327</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>48.5,-60</position>
<output>
<ID>A_equal_B</ID>348 </output>
<output>
<ID>A_greater_B</ID>349 </output>
<output>
<ID>A_less_B</ID>347 </output>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>12 </input>
<input>
<ID>IN_B_0</ID>130 </input>
<input>
<ID>IN_B_1</ID>131 </input>
<input>
<ID>IN_B_2</ID>132 </input>
<input>
<ID>IN_B_3</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>347</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>36,-69</position>
<input>
<ID>ENABLE_0</ID>350 </input>
<input>
<ID>IN_0</ID>346 </input>
<input>
<ID>IN_1</ID>346 </input>
<input>
<ID>IN_2</ID>346 </input>
<input>
<ID>IN_3</ID>349 </input>
<output>
<ID>OUT_0</ID>177 </output>
<output>
<ID>OUT_1</ID>176 </output>
<output>
<ID>OUT_2</ID>175 </output>
<output>
<ID>OUT_3</ID>174 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>348</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>44.5,-69</position>
<input>
<ID>ENABLE_0</ID>351 </input>
<input>
<ID>IN_0</ID>346 </input>
<input>
<ID>IN_1</ID>346 </input>
<input>
<ID>IN_2</ID>346 </input>
<input>
<ID>IN_3</ID>348 </input>
<output>
<ID>OUT_0</ID>177 </output>
<output>
<ID>OUT_1</ID>176 </output>
<output>
<ID>OUT_2</ID>175 </output>
<output>
<ID>OUT_3</ID>174 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>349</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>53,-69</position>
<input>
<ID>ENABLE_0</ID>352 </input>
<input>
<ID>IN_0</ID>346 </input>
<input>
<ID>IN_1</ID>346 </input>
<input>
<ID>IN_2</ID>346 </input>
<input>
<ID>IN_3</ID>347 </input>
<output>
<ID>OUT_0</ID>177 </output>
<output>
<ID>OUT_1</ID>176 </output>
<output>
<ID>OUT_2</ID>175 </output>
<output>
<ID>OUT_3</ID>174 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>351</ID>
<type>FF_GND</type>
<position>56.5,-65</position>
<output>
<ID>OUT_0</ID>346 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>352</ID>
<type>DA_FROM</type>
<position>40,-88</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID GE2D</lparam></gate>
<gate>
<ID>353</ID>
<type>DA_FROM</type>
<position>48.5,-88</position>
<input>
<ID>IN_0</ID>351 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID EQ2D</lparam></gate>
<gate>
<ID>354</ID>
<type>DA_FROM</type>
<position>58,-88</position>
<input>
<ID>IN_0</ID>352 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID LE2D</lparam></gate>
<gate>
<ID>360</ID>
<type>BI_DECODER_4x16</type>
<position>136.5,3.5</position>
<input>
<ID>ENABLE</ID>308 </input>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<input>
<ID>IN_3</ID>54 </input>
<output>
<ID>OUT_0</ID>391 </output>
<output>
<ID>OUT_1</ID>392 </output>
<output>
<ID>OUT_2</ID>393 </output>
<output>
<ID>OUT_3</ID>394 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>361</ID>
<type>DE_TO</type>
<position>141.5,20.5</position>
<input>
<ID>IN_0</ID>394 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>362</ID>
<type>DE_TO</type>
<position>149,20.5</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID GE</lparam></gate>
<gate>
<ID>363</ID>
<type>DE_TO</type>
<position>146.5,20.5</position>
<input>
<ID>IN_0</ID>392 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID EQ</lparam></gate>
<gate>
<ID>364</ID>
<type>DE_TO</type>
<position>144,20.5</position>
<input>
<ID>IN_0</ID>393 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID LE</lparam></gate>
<gate>
<ID>366</ID>
<type>AE_OR2</type>
<position>193,87.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>397 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>371</ID>
<type>DA_FROM</type>
<position>158.5,106.5</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID GE</lparam></gate>
<gate>
<ID>372</ID>
<type>DA_FROM</type>
<position>155.5,106.5</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID EQ</lparam></gate>
<gate>
<ID>373</ID>
<type>DA_FROM</type>
<position>153,106.5</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID LE</lparam></gate>
<gate>
<ID>374</ID>
<type>DE_TO</type>
<position>232,49.5</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID GE2D</lparam></gate>
<gate>
<ID>375</ID>
<type>DE_TO</type>
<position>232,46</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LE2D</lparam></gate>
<gate>
<ID>376</ID>
<type>DE_TO</type>
<position>232,42</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID EQ2D</lparam></gate>
<gate>
<ID>380</ID>
<type>AE_OR3</type>
<position>178.5,56</position>
<input>
<ID>IN_0</ID>370 </input>
<input>
<ID>IN_1</ID>371 </input>
<input>
<ID>IN_2</ID>372 </input>
<output>
<ID>OUT</ID>375 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-26,17,-25</points>
<intersection>-26 4</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-25,18,-25</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>16.5,-26,17,-26</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-4,149,18.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139.5,-4,149,-4</points>
<connection>
<GID>360</GID>
<name>OUT_0</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,105.5,226.5,108</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226.5,108,229.5,108</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-3,146.5,18.5</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139.5,-3,146.5,-3</points>
<connection>
<GID>360</GID>
<name>OUT_1</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23.5,8,-18.5,8</points>
<connection>
<GID>300</GID>
<name>CLK</name></connection>
<connection>
<GID>3</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-2,144,18.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139.5,-2,144,-2</points>
<connection>
<GID>360</GID>
<name>OUT_2</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-23,18,-23</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-1,141.5,18.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139.5,-1,141.5,-1</points>
<connection>
<GID>360</GID>
<name>OUT_3</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107.5,57,117.5,57</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<connection>
<GID>7</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>123.5,58,137.5,58</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107.5,50,117.5,50</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196,87.5,198.5,87.5</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<connection>
<GID>395</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>123.5,51,137.5,51</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-61.5,-2.5,-60</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-60,4.5,-60</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-2.5 0</intersection>
<intersection>4.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>4.5,-61.5,4.5,-50.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-60 1</intersection>
<intersection>-50.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4.5,-50.5,46.5,-50.5</points>
<intersection>4.5 3</intersection>
<intersection>7 9</intersection>
<intersection>21 6</intersection>
<intersection>46.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>21,-56,21,-50.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-50.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>46.5,-56,46.5,-50.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>-50.5 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>7,-50.5,7,-46.5</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>-50.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-61.5,-1.5,-59</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-59,5.5,-59</points>
<connection>
<GID>26</GID>
<name>OUT_1</name></connection>
<intersection>-1.5 0</intersection>
<intersection>5.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>5.5,-61.5,5.5,-51.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>-59 1</intersection>
<intersection>-51.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>5.5,-51.5,45.5,-51.5</points>
<intersection>5.5 3</intersection>
<intersection>20 6</intersection>
<intersection>45.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>20,-56,20,-51.5</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>-51.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>45.5,-56,45.5,-51.5</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>-51.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-61.5,-0.5,-58</points>
<connection>
<GID>28</GID>
<name>IN_2</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-58,6.5,-58</points>
<connection>
<GID>26</GID>
<name>OUT_2</name></connection>
<intersection>-0.5 0</intersection>
<intersection>6.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>6.5,-61.5,6.5,-52.5</points>
<connection>
<GID>47</GID>
<name>IN_2</name></connection>
<intersection>-58 1</intersection>
<intersection>-52.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-52.5,44.5,-52.5</points>
<intersection>6.5 3</intersection>
<intersection>19 6</intersection>
<intersection>44.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>19,-56,19,-52.5</points>
<connection>
<GID>140</GID>
<name>IN_2</name></connection>
<intersection>-52.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>44.5,-56,44.5,-52.5</points>
<connection>
<GID>327</GID>
<name>IN_2</name></connection>
<intersection>-52.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,92,181,103.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181,92,210,92</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-61.5,0.5,-57</points>
<connection>
<GID>28</GID>
<name>IN_3</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-57,7.5,-57</points>
<connection>
<GID>26</GID>
<name>OUT_3</name></connection>
<intersection>0.5 0</intersection>
<intersection>7.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7.5,-61.5,7.5,-53.5</points>
<connection>
<GID>47</GID>
<name>IN_3</name></connection>
<intersection>-57 1</intersection>
<intersection>-53.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>7.5,-53.5,43.5,-53.5</points>
<intersection>7.5 3</intersection>
<intersection>18 7</intersection>
<intersection>43.5 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>18,-56,18,-53.5</points>
<connection>
<GID>140</GID>
<name>IN_3</name></connection>
<intersection>-53.5 6</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>43.5,-56,43.5,-53.5</points>
<connection>
<GID>327</GID>
<name>IN_3</name></connection>
<intersection>-53.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,86.5,207,86.5</points>
<connection>
<GID>395</GID>
<name>OUT</name></connection>
<intersection>207 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>207,86.5,207,90</points>
<intersection>86.5 1</intersection>
<intersection>90 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>207,90,210,90</points>
<connection>
<GID>400</GID>
<name>IN_1</name></connection>
<intersection>207 3</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-24,26,-23</points>
<intersection>-24 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-23,27.5,-23</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-24,26,-24</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-63.5,2.5,-57</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2,-63.5,2.5,-63.5</points>
<connection>
<GID>28</GID>
<name>ENABLE_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-21,26,-19.5</points>
<intersection>-21 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-21,27.5,-21</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-19.5,26,-19.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149.5,36,230,36</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>149.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>149.5,36,149.5,105</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>36 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>226.5,90,229.5,90</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-11,-34.5,-9.5</points>
<intersection>-11 4</intersection>
<intersection>-9.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-36,-11,-34.5,-11</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>-34.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-34.5,-9.5,-33.5,-9.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<intersection>-34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,91,220.5,91</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<connection>
<GID>400</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36,-7.5,-33.5,-7.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<connection>
<GID>405</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107.5,43.5,117.5,43.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,-54,-9,-51</points>
<connection>
<GID>26</GID>
<name>load</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-104.5,34,-104.5</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>32 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>32,-104.5,32,-100.5</points>
<intersection>-104.5 1</intersection>
<intersection>-100.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>28,-100.5,32,-100.5</points>
<connection>
<GID>22</GID>
<name>write_enable</name></connection>
<intersection>32 7</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-96.5,-0.5,-93</points>
<connection>
<GID>64</GID>
<name>load</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-109.5,29.5,-101.5</points>
<intersection>-109.5 1</intersection>
<intersection>-101.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-109.5,34,-109.5</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-101.5,29.5,-101.5</points>
<connection>
<GID>22</GID>
<name>ENABLE_0</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-33.5,223,-33.5</points>
<connection>
<GID>43</GID>
<name>N_in1</name></connection>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<intersection>78 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>78,-33.5,78,-24</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-34.5,223,-34.5</points>
<connection>
<GID>44</GID>
<name>N_in1</name></connection>
<connection>
<GID>40</GID>
<name>N_in0</name></connection>
<intersection>79 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>79,-34.5,79,-24</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-35.5,223,-35.5</points>
<connection>
<GID>45</GID>
<name>N_in1</name></connection>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<intersection>80 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>80,-35.5,80,-24</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-36.5,223,-36.5</points>
<connection>
<GID>46</GID>
<name>N_in1</name></connection>
<connection>
<GID>42</GID>
<name>N_in0</name></connection>
<intersection>81 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>81,-36.5,81,-24</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>123.5,44.5,137.5,44.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>51</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,97.5,116.5,97.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>122.5,98.5,136.5,98.5</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,84.5,116.5,84.5</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9,-63.5,10,-63.5</points>
<connection>
<GID>47</GID>
<name>ENABLE_0</name></connection>
<intersection>10 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>10,-63.5,10,-62</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-63.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-5.5,54,-1</points>
<connection>
<GID>24</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-5.5,61.5,-5.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>34 3</intersection>
<intersection>54 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-5.5,34,6.5</points>
<intersection>-5.5 1</intersection>
<intersection>6.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>34,6.5,39,6.5</points>
<connection>
<GID>54</GID>
<name>IN_4</name></connection>
<intersection>34 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-4.5,53,-1</points>
<connection>
<GID>24</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-4.5,61.5,-4.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>33 3</intersection>
<intersection>53 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,-4.5,33,7.5</points>
<intersection>-4.5 1</intersection>
<intersection>7.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33,7.5,39,7.5</points>
<connection>
<GID>54</GID>
<name>IN_5</name></connection>
<intersection>33 3</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-3.5,52,-1</points>
<connection>
<GID>24</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-3.5,61.5,-3.5</points>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<intersection>32 3</intersection>
<intersection>52 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-3.5,32,8.5</points>
<intersection>-3.5 1</intersection>
<intersection>8.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>32,8.5,39,8.5</points>
<connection>
<GID>54</GID>
<name>IN_6</name></connection>
<intersection>32 3</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-102.5,13,-96.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-102.5,18,-102.5</points>
<connection>
<GID>22</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-18.5,58,-1</points>
<connection>
<GID>24</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-18.5 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-18.5,61.5,-18.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-6.5,58,-6.5</points>
<intersection>38 3</intersection>
<intersection>58 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-6.5,38,2.5</points>
<intersection>-6.5 2</intersection>
<intersection>2.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>38,2.5,39,2.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-17.5,57,-1</points>
<connection>
<GID>24</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-17.5 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-17.5,61.5,-17.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-7.5,57,-7.5</points>
<intersection>37 3</intersection>
<intersection>57 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37,-7.5,37,3.5</points>
<intersection>-7.5 2</intersection>
<intersection>3.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37,3.5,39,3.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>37 3</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-16.5,56,-1</points>
<connection>
<GID>24</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-16.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-16.5,61.5,-16.5</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-8.5,56,-8.5</points>
<intersection>36 3</intersection>
<intersection>56 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-8.5,36,4.5</points>
<intersection>-8.5 2</intersection>
<intersection>4.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,4.5,39,4.5</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>36 3</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-15.5,55,-1</points>
<connection>
<GID>24</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-15.5 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-15.5,61.5,-15.5</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-9.5,55,-9.5</points>
<intersection>35 3</intersection>
<intersection>55 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35,-9.5,35,5.5</points>
<intersection>-9.5 2</intersection>
<intersection>5.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>35,5.5,39,5.5</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<intersection>35 3</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,9.5,49.5,9.5</points>
<connection>
<GID>24</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>54</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,8.5,49.5,8.5</points>
<connection>
<GID>24</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>54</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,7.5,49.5,7.5</points>
<connection>
<GID>24</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>54</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,6.5,49.5,6.5</points>
<connection>
<GID>24</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>54</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,5.5,49.5,5.5</points>
<connection>
<GID>24</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>54</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,4.5,49.5,4.5</points>
<connection>
<GID>24</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>54</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,3.5,49.5,3.5</points>
<connection>
<GID>24</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>54</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,2.5,49.5,2.5</points>
<connection>
<GID>24</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-12,60.5,15.5</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<intersection>-12 4</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,5.5,64.5,5.5</points>
<connection>
<GID>24</GID>
<name>ENABLE_0</name></connection>
<intersection>60.5 0</intersection>
<intersection>64.5 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>60.5,-12,64.5,-12</points>
<intersection>60.5 0</intersection>
<intersection>64.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>64.5,0.5,64.5,5.5</points>
<connection>
<GID>50</GID>
<name>load</name></connection>
<intersection>5.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>64.5,-12.5,64.5,-12</points>
<connection>
<GID>52</GID>
<name>load</name></connection>
<intersection>-12 4</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-20,71,-18.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-18.5,151.5,-18.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection>
<intersection>78 3</intersection>
<intersection>91 13</intersection>
<intersection>131.5 11</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>78,-20,78,-18.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>131.5,-18.5,131.5,-4</points>
<intersection>-18.5 1</intersection>
<intersection>-4 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>131.5,-4,133.5,-4</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>131.5 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>91,-20,91,-18.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-20,72,-17.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-17.5,151.5,-17.5</points>
<connection>
<GID>52</GID>
<name>OUT_1</name></connection>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection>
<intersection>79 3</intersection>
<intersection>90 13</intersection>
<intersection>130.5 11</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>79,-20,79,-17.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>130.5,-17.5,130.5,-3</points>
<intersection>-17.5 1</intersection>
<intersection>-3 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>130.5,-3,133.5,-3</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>130.5 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>90,-22,90,-17.5</points>
<intersection>-22 14</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>90,-22,91,-22</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>90 13</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-20,73,-16.5</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-16.5,151.5,-16.5</points>
<connection>
<GID>52</GID>
<name>OUT_2</name></connection>
<connection>
<GID>67</GID>
<name>IN_2</name></connection>
<intersection>73 0</intersection>
<intersection>80 3</intersection>
<intersection>89 13</intersection>
<intersection>129.5 11</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80,-20,80,-16.5</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>129.5,-16.5,129.5,-2</points>
<intersection>-16.5 1</intersection>
<intersection>-2 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>129.5,-2,133.5,-2</points>
<connection>
<GID>360</GID>
<name>IN_2</name></connection>
<intersection>129.5 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>89,-24,89,-16.5</points>
<intersection>-24 14</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>89,-24,91,-24</points>
<connection>
<GID>100</GID>
<name>IN_2</name></connection>
<intersection>89 13</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-20,74,-15.5</points>
<connection>
<GID>57</GID>
<name>IN_3</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-15.5,128.5,-15.5</points>
<connection>
<GID>52</GID>
<name>OUT_3</name></connection>
<intersection>74 0</intersection>
<intersection>81 3</intersection>
<intersection>88 11</intersection>
<intersection>128.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>81,-20,81,-15.5</points>
<connection>
<GID>59</GID>
<name>IN_3</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>128.5,-15.5,128.5,-1</points>
<intersection>-15.5 1</intersection>
<intersection>-1 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>128.5,-1,133.5,-1</points>
<connection>
<GID>360</GID>
<name>IN_3</name></connection>
<intersection>128.5 8</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>88,-26,88,-15.5</points>
<intersection>-26 12</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>88,-26,91,-26</points>
<connection>
<GID>100</GID>
<name>IN_3</name></connection>
<intersection>88 11</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-22,76.5,-14.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-22,76.5,-22</points>
<connection>
<GID>57</GID>
<name>ENABLE_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-22,84.5,-14.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-22,84.5,-22</points>
<connection>
<GID>59</GID>
<name>ENABLE_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,-2.5,101,-2.5</points>
<connection>
<GID>50</GID>
<name>OUT_3</name></connection>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>95 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>95,-2.5,95,15.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-2.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,-3.5,101,-3.5</points>
<connection>
<GID>50</GID>
<name>OUT_2</name></connection>
<connection>
<GID>62</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,-4.5,101,-4.5</points>
<connection>
<GID>50</GID>
<name>OUT_1</name></connection>
<connection>
<GID>62</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,-5.5,101,-5.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<connection>
<GID>62</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-101.5,14,-96.5</points>
<connection>
<GID>76</GID>
<name>OUT_1</name></connection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-101.5,18,-101.5</points>
<connection>
<GID>22</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>86</GID>
<name>OUT_1</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-100.5,15,-96.5</points>
<connection>
<GID>76</GID>
<name>OUT_2</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-100.5,18,-100.5</points>
<connection>
<GID>22</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>86</GID>
<name>OUT_2</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-99.5,16,-96.5</points>
<connection>
<GID>76</GID>
<name>OUT_3</name></connection>
<intersection>-99.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-99.5,18,-99.5</points>
<connection>
<GID>22</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>86</GID>
<name>OUT_3</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-99.5,5.5,-99.5</points>
<connection>
<GID>86</GID>
<name>IN_3</name></connection>
<connection>
<GID>64</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-100.5,5.5,-100.5</points>
<connection>
<GID>86</GID>
<name>IN_2</name></connection>
<connection>
<GID>64</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-101.5,5.5,-101.5</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-102.5,5.5,-102.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-23,99,-23</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>100</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>167,72.5,229.5,72.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>167 3</intersection>
<intersection>218.5 17</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>167,72.5,167,104</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>72.5 1</intersection>
<intersection>75 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>167,75,192,75</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>167 3</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>218.5,72.5,218.5,89</points>
<intersection>72.5 1</intersection>
<intersection>89 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>218.5,89,220.5,89</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>218.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>198,76,229.5,76</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173.5,95,229.5,95</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>173.5 20</intersection>
<intersection>190 25</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>173.5,95,173.5,103.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>95 1</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>190,88.5,190,95</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>95 1</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>170,77,170,103.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>77 23</intersection>
<intersection>83.5 12</intersection>
<intersection>98 36</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>170,83.5,229.5,83.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>170 9</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>170,77,192,77</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>170 9</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>170,98,188,98</points>
<connection>
<GID>261</GID>
<name>IN_1</name></connection>
<intersection>170 9</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,0,-13,9.5</points>
<connection>
<GID>23</GID>
<name>clock</name></connection>
<intersection>0 2</intersection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,8,-13,8</points>
<connection>
<GID>3</GID>
<name>N_in1</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13,0,-12,0</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>122.5,85.5,136.5,85.5</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<connection>
<GID>90</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-98,7.5,-90</points>
<connection>
<GID>86</GID>
<name>ENABLE_0</name></connection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-90,24,-90</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>7.5 0</intersection>
<intersection>22.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>22.5,-94.5,22.5,-90</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-90 1</intersection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,90.5,116.5,90.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-5.5,126.5,18</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-5.5,126.5,-5.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-4.5,124,18</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-4.5,124,-4.5</points>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection>
<intersection>124 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-10.5,121.5,18</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-10.5 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-3.5,121.5,-3.5</points>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-10.5,144,-10.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-12.5,119,18</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-12.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-2.5,119,-2.5</points>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,-12.5,144,-12.5</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-1.5,116.5,18</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-1.5,116.5,-1.5</points>
<connection>
<GID>62</GID>
<name>OUT_4</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-0.5,114,18</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-0.5,114,-0.5</points>
<connection>
<GID>62</GID>
<name>OUT_5</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-94.5,18.5,-94.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<connection>
<GID>76</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,12.5,-7,12.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,13.5,-7,13.5</points>
<connection>
<GID>23</GID>
<name>OUT_1</name></connection>
<connection>
<GID>49</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,14.5,-7,14.5</points>
<connection>
<GID>23</GID>
<name>OUT_2</name></connection>
<connection>
<GID>49</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-26,3.5,7.5,3.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>1 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1,3.5,1,5.5</points>
<intersection>3.5 1</intersection>
<intersection>5.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-3,5.5,1,5.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>1 7</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>122.5,91.5,136.5,91.5</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-11.5,163.5,-5.5</points>
<intersection>-11.5 2</intersection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-5.5,170.5,-5.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-11.5,163.5,-11.5</points>
<connection>
<GID>67</GID>
<name>OUT_7</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-12.5,164.5,-8</points>
<intersection>-12.5 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164.5,-8,170.5,-8</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-12.5,164.5,-12.5</points>
<connection>
<GID>67</GID>
<name>OUT_6</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-11,64.5,-11</points>
<intersection>53 5</intersection>
<intersection>64.5 8</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>53,-21.5,53,-11</points>
<intersection>-21.5 7</intersection>
<intersection>-16 15</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>53,-21.5,64.5,-21.5</points>
<connection>
<GID>52</GID>
<name>clock</name></connection>
<intersection>53 5</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>64.5,-11,64.5,-8.5</points>
<connection>
<GID>50</GID>
<name>clock</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>33.5,-16,53,-16</points>
<intersection>33.5 16</intersection>
<intersection>53 5</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>33.5,-22,33.5,-16</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<intersection>-16 15</intersection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,10,0,12.5</points>
<intersection>10 1</intersection>
<intersection>12.5 12</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,10,7,10</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-1,12.5,0,12.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,6.5,-11,9.5</points>
<connection>
<GID>23</GID>
<name>clear</name></connection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,6.5,-9,6.5</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-22.5,44,0.5</points>
<connection>
<GID>54</GID>
<name>clear</name></connection>
<intersection>-22.5 1</intersection>
<intersection>-10.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-22.5,66.5,-22.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection>
<intersection>66.5 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>44,-10.5,66.5,-10.5</points>
<intersection>44 0</intersection>
<intersection>66.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>66.5,-10.5,66.5,-8.5</points>
<connection>
<GID>50</GID>
<name>clear</name></connection>
<intersection>-10.5 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>66.5,-22.5,66.5,-21.5</points>
<connection>
<GID>52</GID>
<name>clear</name></connection>
<intersection>-22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,18.5,7,18.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>1.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>1.5,7.5,1.5,18.5</points>
<intersection>7.5 9</intersection>
<intersection>15.5 7</intersection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1,15.5,1.5,15.5</points>
<connection>
<GID>49</GID>
<name>OUT_3</name></connection>
<intersection>1.5 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-3,7.5,1.5,7.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>1.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,18.5,-12,21.5</points>
<connection>
<GID>23</GID>
<name>count_enable</name></connection>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<intersection>19.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-12,19.5,-7,19.5</points>
<connection>
<GID>49</GID>
<name>ENABLE</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-27.5,71,-24</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17.5,-27.5,223,-27.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>15</GID>
<name>N_in1</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-28.5,72,-24</points>
<connection>
<GID>57</GID>
<name>OUT_1</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17.5,-28.5,223,-28.5</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<connection>
<GID>16</GID>
<name>N_in1</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-29.5,73,-24</points>
<connection>
<GID>57</GID>
<name>OUT_2</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17.5,-29.5,223,-29.5</points>
<connection>
<GID>11</GID>
<name>N_in0</name></connection>
<connection>
<GID>17</GID>
<name>N_in1</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164,-23.5,164,-18.5</points>
<intersection>-23.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164,-23.5,170,-23.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>164 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-18.5,164,-18.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>164 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-21,165,-17.5</points>
<intersection>-21 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-21,170,-21</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-17.5,165,-17.5</points>
<connection>
<GID>67</GID>
<name>OUT_1</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-18.5,166,-16.5</points>
<intersection>-18.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-18.5,170,-18.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-16.5,166,-16.5</points>
<connection>
<GID>67</GID>
<name>OUT_2</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,-15.5,170,-15.5</points>
<connection>
<GID>67</GID>
<name>OUT_3</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-30.5,74,-24</points>
<connection>
<GID>57</GID>
<name>OUT_3</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17.5,-30.5,223,-30.5</points>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<connection>
<GID>18</GID>
<name>N_in1</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-61.5,74.5,-48.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-60 1</intersection>
<intersection>-48.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-60,74.5,-60</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28,-48.5,74.5,-48.5</points>
<intersection>28 4</intersection>
<intersection>53.5 5</intersection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>28,-56,28,-48.5</points>
<connection>
<GID>140</GID>
<name>IN_B_0</name></connection>
<intersection>-48.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>53.5,-56,53.5,-48.5</points>
<connection>
<GID>327</GID>
<name>IN_B_0</name></connection>
<intersection>-48.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-61.5,75.5,-47.5</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>-59 1</intersection>
<intersection>-47.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-59,75.5,-59</points>
<connection>
<GID>130</GID>
<name>OUT_1</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-47.5,75.5,-47.5</points>
<intersection>27 4</intersection>
<intersection>52.5 5</intersection>
<intersection>75.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27,-56,27,-47.5</points>
<connection>
<GID>140</GID>
<name>IN_B_1</name></connection>
<intersection>-47.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>52.5,-56,52.5,-47.5</points>
<connection>
<GID>327</GID>
<name>IN_B_1</name></connection>
<intersection>-47.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-61.5,76.5,-46.5</points>
<connection>
<GID>131</GID>
<name>IN_2</name></connection>
<intersection>-58 1</intersection>
<intersection>-46.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-58,76.5,-58</points>
<connection>
<GID>130</GID>
<name>OUT_2</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-46.5,76.5,-46.5</points>
<intersection>26 4</intersection>
<intersection>51.5 5</intersection>
<intersection>76.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>26,-56,26,-46.5</points>
<connection>
<GID>140</GID>
<name>IN_B_2</name></connection>
<intersection>-46.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>51.5,-56,51.5,-46.5</points>
<connection>
<GID>327</GID>
<name>IN_B_2</name></connection>
<intersection>-46.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-61.5,77.5,-45.5</points>
<connection>
<GID>131</GID>
<name>IN_3</name></connection>
<intersection>-57 1</intersection>
<intersection>-45.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-57,77.5,-57</points>
<connection>
<GID>130</GID>
<name>OUT_3</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25,-45.5,77.5,-45.5</points>
<intersection>25 4</intersection>
<intersection>50.5 5</intersection>
<intersection>77.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>25,-56,25,-45.5</points>
<connection>
<GID>140</GID>
<name>IN_B_3</name></connection>
<intersection>-45.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>50.5,-56,50.5,-45.5</points>
<connection>
<GID>327</GID>
<name>IN_B_3</name></connection>
<intersection>-45.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-63.5,79.5,-57</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>79,-63.5,79.5,-63.5</points>
<connection>
<GID>131</GID>
<name>ENABLE_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-62.5,63.5,-60</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-60,65,-60</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-62.5,62.5,-59</points>
<connection>
<GID>133</GID>
<name>OUT_1</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-59,65,-59</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-62.5,61.5,-58</points>
<connection>
<GID>133</GID>
<name>OUT_2</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-58,65,-58</points>
<connection>
<GID>130</GID>
<name>IN_2</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-62.5,60.5,-57</points>
<connection>
<GID>133</GID>
<name>OUT_3</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-57,65,-57</points>
<connection>
<GID>130</GID>
<name>IN_3</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-64.5,58,-62</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-64.5,59,-64.5</points>
<connection>
<GID>133</GID>
<name>ENABLE_0</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-80.5,205,-80.5</points>
<connection>
<GID>200</GID>
<name>N_in0</name></connection>
<connection>
<GID>165</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-54,68,-52.5</points>
<connection>
<GID>130</GID>
<name>load</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,-52.5,68,-52.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-65.5,21.5,-64</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<connection>
<GID>140</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-65.5,22.5,-64</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<connection>
<GID>140</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-65.5,23.5,-64</points>
<connection>
<GID>141</GID>
<name>IN_2</name></connection>
<connection>
<GID>140</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-65.5,24.5,-64</points>
<connection>
<GID>141</GID>
<name>IN_3</name></connection>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-67.5,32.5,-65.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-67.5,32.5,-67.5</points>
<connection>
<GID>141</GID>
<name>ENABLE_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-81.5,205,-81.5</points>
<connection>
<GID>201</GID>
<name>N_in0</name></connection>
<connection>
<GID>166</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-82.5,205,-82.5</points>
<connection>
<GID>202</GID>
<name>N_in0</name></connection>
<connection>
<GID>167</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-41,223,-41</points>
<connection>
<GID>145</GID>
<name>N_in0</name></connection>
<connection>
<GID>147</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-40,223,-40</points>
<connection>
<GID>144</GID>
<name>N_in0</name></connection>
<connection>
<GID>146</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-107,42.5,-107</points>
<intersection>-0.5 22</intersection>
<intersection>42.5 23</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-0.5,-107,-0.5,-105.5</points>
<connection>
<GID>64</GID>
<name>clock</name></connection>
<intersection>-107 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>42.5,-107,42.5,-99.5</points>
<intersection>-107 1</intersection>
<intersection>-99.5 25</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>28,-99.5,43.5,-99.5</points>
<connection>
<GID>22</GID>
<name>write_clock</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>42.5 23</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150,-11.5,151.5,-11.5</points>
<connection>
<GID>67</GID>
<name>ENABLE</name></connection>
<connection>
<GID>152</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-27.5,225,-21</points>
<connection>
<GID>8</GID>
<name>N_in1</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-21,229.5,-21</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,-28.5,226,-23.5</points>
<intersection>-28.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,-23.5,229.5,-23.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225,-28.5,226,-28.5</points>
<connection>
<GID>10</GID>
<name>N_in1</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-29.5,227,-26</points>
<intersection>-29.5 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,-26,229.5,-26</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>227 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225,-29.5,227,-29.5</points>
<connection>
<GID>11</GID>
<name>N_in1</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>229.5,-30.5,229.5,-28.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-30.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>225,-30.5,229.5,-30.5</points>
<connection>
<GID>12</GID>
<name>N_in1</name></connection>
<intersection>229.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-33.5,227,-31.5</points>
<intersection>-33.5 2</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>225,-33.5,227,-33.5</points>
<connection>
<GID>39</GID>
<name>N_in1</name></connection>
<intersection>227 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>227,-31.5,229.5,-31.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-34.5,229.5,-34.5</points>
<connection>
<GID>40</GID>
<name>N_in1</name></connection>
<intersection>229.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,-34.5,229.5,-34</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,-36.5,226,-35.5</points>
<intersection>-36.5 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,-36.5,229.5,-36.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225,-35.5,226,-35.5</points>
<connection>
<GID>41</GID>
<name>N_in1</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,-39,226,-36.5</points>
<intersection>-39 1</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,-39,229.5,-39</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225,-36.5,226,-36.5</points>
<connection>
<GID>42</GID>
<name>N_in1</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-43.5,227,-40</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>225,-40,227,-40</points>
<connection>
<GID>144</GID>
<name>N_in1</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,-47,226,-41</points>
<intersection>-47 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,-47,227,-47</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225,-41,226,-41</points>
<connection>
<GID>145</GID>
<name>N_in1</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-83.5,205,-83.5</points>
<connection>
<GID>203</GID>
<name>N_in0</name></connection>
<connection>
<GID>168</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,-77.5,-25,-30.5</points>
<intersection>-77.5 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-77.5,-22,-77.5</points>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-25,-30.5,-19.5,-30.5</points>
<connection>
<GID>18</GID>
<name>N_in0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26,-76.5,-26,-29.5</points>
<intersection>-76.5 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26,-76.5,-22,-76.5</points>
<connection>
<GID>139</GID>
<name>N_in0</name></connection>
<intersection>-26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26,-29.5,-19.5,-29.5</points>
<connection>
<GID>17</GID>
<name>N_in0</name></connection>
<intersection>-26 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,-75.5,-27,-28.5</points>
<intersection>-75.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27,-75.5,-22,-75.5</points>
<connection>
<GID>136</GID>
<name>N_in0</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27,-28.5,-19.5,-28.5</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<intersection>-27 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-74.5,-28,-27.5</points>
<intersection>-74.5 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28,-74.5,-22,-74.5</points>
<connection>
<GID>135</GID>
<name>N_in0</name></connection>
<intersection>-28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,-27.5,-19.5,-27.5</points>
<connection>
<GID>15</GID>
<name>N_in0</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30.5,-83.5,-30.5,-36.5</points>
<intersection>-83.5 1</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30.5,-83.5,-22,-83.5</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<intersection>-30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-30.5,-36.5,-19.5,-36.5</points>
<connection>
<GID>46</GID>
<name>N_in0</name></connection>
<intersection>-30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31.5,-82.5,-31.5,-35.5</points>
<intersection>-82.5 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-31.5,-82.5,-22,-82.5</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<intersection>-31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-31.5,-35.5,-19.5,-35.5</points>
<connection>
<GID>45</GID>
<name>N_in0</name></connection>
<intersection>-31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-81.5,-32.5,-34.5</points>
<intersection>-81.5 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,-81.5,-22,-81.5</points>
<connection>
<GID>153</GID>
<name>N_in0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-32.5,-34.5,-19.5,-34.5</points>
<connection>
<GID>44</GID>
<name>N_in0</name></connection>
<intersection>-32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-80.5,-33.5,-33.5</points>
<intersection>-80.5 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,-80.5,-22,-80.5</points>
<connection>
<GID>151</GID>
<name>N_in0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,-33.5,-19.5,-33.5</points>
<connection>
<GID>43</GID>
<name>N_in0</name></connection>
<intersection>-33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-74.5,-13.5,-60</points>
<intersection>-74.5 1</intersection>
<intersection>-60 21</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-74.5,80.5,-74.5</points>
<connection>
<GID>135</GID>
<name>N_in1</name></connection>
<connection>
<GID>157</GID>
<name>N_in0</name></connection>
<intersection>-13.5 0</intersection>
<intersection>-8 16</intersection>
<intersection>-2.5 3</intersection>
<intersection>24.5 4</intersection>
<intersection>37.5 12</intersection>
<intersection>46 14</intersection>
<intersection>54.5 15</intersection>
<intersection>63.5 5</intersection>
<intersection>74.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2.5,-74.5,-2.5,-65.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>24.5,-74.5,24.5,-69.5</points>
<connection>
<GID>141</GID>
<name>OUT_3</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>63.5,-74.5,63.5,-66.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>74.5,-74.5,74.5,-65.5</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>37.5,-74.5,37.5,-71</points>
<connection>
<GID>347</GID>
<name>OUT_3</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>46,-74.5,46,-71</points>
<connection>
<GID>348</GID>
<name>OUT_3</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>54.5,-74.5,54.5,-71</points>
<connection>
<GID>349</GID>
<name>OUT_3</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-8,-116,-8,-74.5</points>
<intersection>-116 17</intersection>
<intersection>-102.5 22</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-8,-116,24.5,-116</points>
<intersection>-8 16</intersection>
<intersection>24.5 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>24.5,-116,24.5,-106</points>
<connection>
<GID>22</GID>
<name>DATA_IN_0</name></connection>
<connection>
<GID>22</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-116 17</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-13.5,-60,-12,-60</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-8,-102.5,-3.5,-102.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-8 16</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-75.5,-14.5,-59</points>
<intersection>-75.5 1</intersection>
<intersection>-59 20</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-75.5,80.5,-75.5</points>
<connection>
<GID>136</GID>
<name>N_in1</name></connection>
<connection>
<GID>158</GID>
<name>N_in0</name></connection>
<intersection>-14.5 0</intersection>
<intersection>-7 15</intersection>
<intersection>-1.5 2</intersection>
<intersection>23.5 3</intersection>
<intersection>36.5 12</intersection>
<intersection>45 13</intersection>
<intersection>53.5 14</intersection>
<intersection>62.5 4</intersection>
<intersection>75.5 5</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-1.5,-75.5,-1.5,-65.5</points>
<connection>
<GID>28</GID>
<name>OUT_1</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>23.5,-75.5,23.5,-69.5</points>
<connection>
<GID>141</GID>
<name>OUT_2</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>62.5,-75.5,62.5,-66.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>75.5,-75.5,75.5,-65.5</points>
<connection>
<GID>131</GID>
<name>OUT_1</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>36.5,-75.5,36.5,-71</points>
<connection>
<GID>347</GID>
<name>OUT_2</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>45,-75.5,45,-71</points>
<connection>
<GID>348</GID>
<name>OUT_2</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>53.5,-75.5,53.5,-71</points>
<connection>
<GID>349</GID>
<name>OUT_2</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-7,-115,-7,-75.5</points>
<intersection>-115 16</intersection>
<intersection>-101.5 21</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-7,-115,23.5,-115</points>
<intersection>-7 15</intersection>
<intersection>23.5 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>23.5,-115,23.5,-106</points>
<connection>
<GID>22</GID>
<name>DATA_IN_1</name></connection>
<connection>
<GID>22</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-115 16</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-14.5,-59,-12,-59</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-7,-101.5,-3.5,-101.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>-7 15</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-76.5,-15.5,-58</points>
<intersection>-76.5 1</intersection>
<intersection>-58 19</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-76.5,80.5,-76.5</points>
<connection>
<GID>139</GID>
<name>N_in1</name></connection>
<connection>
<GID>159</GID>
<name>N_in0</name></connection>
<intersection>-15.5 0</intersection>
<intersection>-6 14</intersection>
<intersection>-0.5 2</intersection>
<intersection>22.5 3</intersection>
<intersection>35.5 11</intersection>
<intersection>44 12</intersection>
<intersection>52.5 13</intersection>
<intersection>61.5 4</intersection>
<intersection>76.5 5</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-0.5,-76.5,-0.5,-65.5</points>
<connection>
<GID>28</GID>
<name>OUT_2</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-76.5,22.5,-69.5</points>
<connection>
<GID>141</GID>
<name>OUT_1</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>61.5,-76.5,61.5,-66.5</points>
<connection>
<GID>133</GID>
<name>IN_2</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>76.5,-76.5,76.5,-65.5</points>
<connection>
<GID>131</GID>
<name>OUT_2</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>35.5,-76.5,35.5,-71</points>
<connection>
<GID>347</GID>
<name>OUT_1</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>44,-76.5,44,-71</points>
<connection>
<GID>348</GID>
<name>OUT_1</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>52.5,-76.5,52.5,-71</points>
<connection>
<GID>349</GID>
<name>OUT_1</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-6,-114,-6,-76.5</points>
<intersection>-114 15</intersection>
<intersection>-100.5 20</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-6,-114,22.5,-114</points>
<intersection>-6 14</intersection>
<intersection>22.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>22.5,-114,22.5,-106</points>
<connection>
<GID>22</GID>
<name>DATA_IN_2</name></connection>
<connection>
<GID>22</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-114 15</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-15.5,-58,-12,-58</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-6,-100.5,-3.5,-100.5</points>
<connection>
<GID>64</GID>
<name>IN_2</name></connection>
<intersection>-6 14</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-77.5,-16.5,-57</points>
<intersection>-77.5 1</intersection>
<intersection>-57 20</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-77.5,80.5,-77.5</points>
<connection>
<GID>148</GID>
<name>N_in1</name></connection>
<connection>
<GID>160</GID>
<name>N_in0</name></connection>
<intersection>-16.5 0</intersection>
<intersection>-5 16</intersection>
<intersection>0.5 2</intersection>
<intersection>21.5 3</intersection>
<intersection>34.5 13</intersection>
<intersection>43 14</intersection>
<intersection>51.5 15</intersection>
<intersection>60.5 4</intersection>
<intersection>77.5 5</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>0.5,-77.5,0.5,-65.5</points>
<connection>
<GID>28</GID>
<name>OUT_3</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>21.5,-77.5,21.5,-69.5</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>60.5,-77.5,60.5,-66.5</points>
<connection>
<GID>133</GID>
<name>IN_3</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>77.5,-77.5,77.5,-65.5</points>
<connection>
<GID>131</GID>
<name>OUT_3</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>34.5,-77.5,34.5,-71</points>
<connection>
<GID>347</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>43,-77.5,43,-71</points>
<connection>
<GID>348</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>51.5,-77.5,51.5,-71</points>
<connection>
<GID>349</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-5,-113,-5,-77.5</points>
<intersection>-113 17</intersection>
<intersection>-99.5 22</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-5,-113,21.5,-113</points>
<intersection>-5 16</intersection>
<intersection>21.5 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>21.5,-113,21.5,-106</points>
<connection>
<GID>22</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>22</GID>
<name>DATA_IN_3</name></connection>
<intersection>-113 17</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-16.5,-57,-12,-57</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>-16.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-5,-99.5,-3.5,-99.5</points>
<connection>
<GID>64</GID>
<name>IN_3</name></connection>
<intersection>-5 16</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-80.5,4.5,-65.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-80.5,80.5,-80.5</points>
<connection>
<GID>151</GID>
<name>N_in1</name></connection>
<connection>
<GID>165</GID>
<name>N_in0</name></connection>
<intersection>4.5 0</intersection>
<intersection>13 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>13,-92.5,13,-80.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-81.5,5.5,-65.5</points>
<connection>
<GID>47</GID>
<name>OUT_1</name></connection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-81.5,80.5,-81.5</points>
<connection>
<GID>153</GID>
<name>N_in1</name></connection>
<connection>
<GID>166</GID>
<name>N_in0</name></connection>
<intersection>5.5 0</intersection>
<intersection>14 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>14,-92.5,14,-81.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-81.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-82.5,6.5,-65.5</points>
<connection>
<GID>47</GID>
<name>OUT_2</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-82.5,80.5,-82.5</points>
<connection>
<GID>154</GID>
<name>N_in1</name></connection>
<connection>
<GID>167</GID>
<name>N_in0</name></connection>
<intersection>6.5 0</intersection>
<intersection>15 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>15,-92.5,15,-82.5</points>
<connection>
<GID>76</GID>
<name>IN_2</name></connection>
<intersection>-82.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-83.5,7.5,-65.5</points>
<connection>
<GID>47</GID>
<name>OUT_3</name></connection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-83.5,80.5,-83.5</points>
<connection>
<GID>155</GID>
<name>N_in1</name></connection>
<connection>
<GID>168</GID>
<name>N_in0</name></connection>
<intersection>7.5 0</intersection>
<intersection>16 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>16,-92.5,16,-83.5</points>
<connection>
<GID>76</GID>
<name>IN_3</name></connection>
<intersection>-83.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,62,230,62</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>161.5 12</intersection>
<intersection>187 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>187,62,187,86.5</points>
<intersection>62 1</intersection>
<intersection>86.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>187,86.5,190,86.5</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>187 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>161.5,62,161.5,104</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>62 1</intersection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>122.5,112,136,112</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,86.5,111,115</points>
<intersection>86.5 9</intersection>
<intersection>92.5 10</intersection>
<intersection>99.5 6</intersection>
<intersection>105.5 4</intersection>
<intersection>113 1</intersection>
<intersection>115 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,113,116.5,113</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,115,111,115</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,105.5,116.5,105.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>111,99.5,116.5,99.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>111,86.5,116.5,86.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111,92.5,116.5,92.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,110,114,111</points>
<intersection>110 2</intersection>
<intersection>111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,111,116.5,111</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>114 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106,110,114,110</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-72,68,-63</points>
<connection>
<GID>130</GID>
<name>clock</name></connection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9,-72,199,-72</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>-9 3</intersection>
<intersection>68 0</intersection>
<intersection>103.5 12</intersection>
<intersection>130.5 11</intersection>
<intersection>157.5 10</intersection>
<intersection>186 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-9,-72,-9,-63</points>
<connection>
<GID>26</GID>
<name>clock</name></connection>
<intersection>-72 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>186,-72,186,-63</points>
<connection>
<GID>181</GID>
<name>clock</name></connection>
<intersection>-72 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>157.5,-72,157.5,-62.5</points>
<connection>
<GID>209</GID>
<name>clock</name></connection>
<intersection>-72 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>130.5,-72,130.5,-62</points>
<connection>
<GID>216</GID>
<name>clock</name></connection>
<intersection>-72 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>103.5,-72,103.5,-62</points>
<connection>
<GID>223</GID>
<name>clock</name></connection>
<intersection>-72 1</intersection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,-61.5,192.5,-60</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-60,192.5,-60</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<intersection>192.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,-61.5,193.5,-59</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-59,193.5,-59</points>
<connection>
<GID>181</GID>
<name>OUT_1</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-61.5,194.5,-58</points>
<connection>
<GID>182</GID>
<name>IN_2</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-58,194.5,-58</points>
<connection>
<GID>181</GID>
<name>OUT_2</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-61.5,195.5,-57</points>
<connection>
<GID>182</GID>
<name>IN_3</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-57,195.5,-57</points>
<connection>
<GID>181</GID>
<name>OUT_3</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-63.5,197.5,-57</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>197,-63.5,197.5,-63.5</points>
<connection>
<GID>182</GID>
<name>ENABLE_0</name></connection>
<intersection>197.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>181.5,-54,186,-54</points>
<connection>
<GID>181</GID>
<name>load</name></connection>
<intersection>181.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>181.5,-54,181.5,-51.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-74.5,205,-74.5</points>
<connection>
<GID>192</GID>
<name>N_in0</name></connection>
<connection>
<GID>157</GID>
<name>N_in1</name></connection>
<intersection>99 10</intersection>
<intersection>110 14</intersection>
<intersection>126 13</intersection>
<intersection>137 12</intersection>
<intersection>153 11</intersection>
<intersection>164 8</intersection>
<intersection>181.5 5</intersection>
<intersection>192.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>181.5,-74.5,181.5,-60</points>
<intersection>-74.5 1</intersection>
<intersection>-60 26</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>192.5,-74.5,192.5,-65.5</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>164,-74.5,164,-65</points>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>99,-74.5,99,-59</points>
<intersection>-74.5 1</intersection>
<intersection>-59 20</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>153,-74.5,153,-59.5</points>
<intersection>-74.5 1</intersection>
<intersection>-59.5 25</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>137,-74.5,137,-64.5</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>126,-74.5,126,-59</points>
<intersection>-74.5 1</intersection>
<intersection>-59 24</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>110,-74.5,110,-64.5</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>99,-59,100.5,-59</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>99 10</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>126,-59,127.5,-59</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>126 13</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>153,-59.5,154.5,-59.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>153 11</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>181.5,-60,183,-60</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>181.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-75.5,205,-75.5</points>
<connection>
<GID>193</GID>
<name>N_in0</name></connection>
<connection>
<GID>158</GID>
<name>N_in1</name></connection>
<intersection>98 9</intersection>
<intersection>111 13</intersection>
<intersection>125 12</intersection>
<intersection>138 11</intersection>
<intersection>152 10</intersection>
<intersection>165 7</intersection>
<intersection>180.5 4</intersection>
<intersection>193.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>180.5,-75.5,180.5,-59</points>
<intersection>-75.5 1</intersection>
<intersection>-59 21</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>193.5,-75.5,193.5,-65.5</points>
<connection>
<GID>182</GID>
<name>OUT_1</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>165,-75.5,165,-65</points>
<connection>
<GID>210</GID>
<name>OUT_1</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>98,-75.5,98,-58</points>
<intersection>-75.5 1</intersection>
<intersection>-58 18</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>152,-75.5,152,-58.5</points>
<intersection>-75.5 1</intersection>
<intersection>-58.5 20</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>138,-75.5,138,-64.5</points>
<connection>
<GID>217</GID>
<name>OUT_1</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>125,-75.5,125,-58</points>
<intersection>-75.5 1</intersection>
<intersection>-58 19</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>111,-75.5,111,-64.5</points>
<connection>
<GID>224</GID>
<name>OUT_1</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>98,-58,100.5,-58</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<intersection>98 9</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>125,-58,127.5,-58</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>125 12</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>152,-58.5,154.5,-58.5</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>152 10</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>180.5,-59,183,-59</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>180.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-76.5,205,-76.5</points>
<connection>
<GID>194</GID>
<name>N_in0</name></connection>
<connection>
<GID>159</GID>
<name>N_in1</name></connection>
<intersection>97 9</intersection>
<intersection>112 13</intersection>
<intersection>124 12</intersection>
<intersection>139 11</intersection>
<intersection>151 10</intersection>
<intersection>166 7</intersection>
<intersection>179.5 4</intersection>
<intersection>194.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>179.5,-76.5,179.5,-58</points>
<intersection>-76.5 1</intersection>
<intersection>-58 21</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>194.5,-76.5,194.5,-65.5</points>
<connection>
<GID>182</GID>
<name>OUT_2</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>166,-76.5,166,-65</points>
<connection>
<GID>210</GID>
<name>OUT_2</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>97,-76.5,97,-57</points>
<intersection>-76.5 1</intersection>
<intersection>-57 18</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>151,-76.5,151,-57.5</points>
<intersection>-76.5 1</intersection>
<intersection>-57.5 20</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>139,-76.5,139,-64.5</points>
<connection>
<GID>217</GID>
<name>OUT_2</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>124,-76.5,124,-57</points>
<intersection>-76.5 1</intersection>
<intersection>-57 19</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>112,-76.5,112,-64.5</points>
<connection>
<GID>224</GID>
<name>OUT_2</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>97,-57,100.5,-57</points>
<connection>
<GID>223</GID>
<name>IN_2</name></connection>
<intersection>97 9</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>124,-57,127.5,-57</points>
<connection>
<GID>216</GID>
<name>IN_2</name></connection>
<intersection>124 12</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>151,-57.5,154.5,-57.5</points>
<connection>
<GID>209</GID>
<name>IN_2</name></connection>
<intersection>151 10</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>179.5,-58,183,-58</points>
<connection>
<GID>181</GID>
<name>IN_2</name></connection>
<intersection>179.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-77.5,205,-77.5</points>
<connection>
<GID>195</GID>
<name>N_in0</name></connection>
<connection>
<GID>160</GID>
<name>N_in1</name></connection>
<intersection>96 9</intersection>
<intersection>113 16</intersection>
<intersection>123 14</intersection>
<intersection>140 13</intersection>
<intersection>150 10</intersection>
<intersection>167 7</intersection>
<intersection>178.5 4</intersection>
<intersection>195.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>178.5,-77.5,178.5,-57</points>
<intersection>-77.5 1</intersection>
<intersection>-57 27</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>195.5,-77.5,195.5,-65.5</points>
<connection>
<GID>182</GID>
<name>OUT_3</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>167,-77.5,167,-65</points>
<connection>
<GID>210</GID>
<name>OUT_3</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>96,-77.5,96,-56</points>
<intersection>-77.5 1</intersection>
<intersection>-56 24</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>150,-77.5,150,-56.5</points>
<intersection>-77.5 1</intersection>
<intersection>-56.5 26</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>140,-77.5,140,-64.5</points>
<connection>
<GID>217</GID>
<name>OUT_3</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>123,-77.5,123,-56</points>
<intersection>-77.5 1</intersection>
<intersection>-56 25</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>113,-77.5,113,-64.5</points>
<connection>
<GID>224</GID>
<name>OUT_3</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>96,-56,100.5,-56</points>
<connection>
<GID>223</GID>
<name>IN_3</name></connection>
<intersection>96 9</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>123,-56,127.5,-56</points>
<connection>
<GID>216</GID>
<name>IN_3</name></connection>
<intersection>123 14</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>150,-56.5,154.5,-56.5</points>
<connection>
<GID>209</GID>
<name>IN_3</name></connection>
<intersection>150 10</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>178.5,-57,183,-57</points>
<connection>
<GID>181</GID>
<name>IN_3</name></connection>
<intersection>178.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164,-61,164,-59.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-59.5,164,-59.5</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>164 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-61,165,-58.5</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-58.5,165,-58.5</points>
<connection>
<GID>209</GID>
<name>OUT_1</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-61,166,-57.5</points>
<connection>
<GID>210</GID>
<name>IN_2</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-57.5,166,-57.5</points>
<connection>
<GID>209</GID>
<name>OUT_2</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-61,167,-56.5</points>
<connection>
<GID>210</GID>
<name>IN_3</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-56.5,167,-56.5</points>
<connection>
<GID>209</GID>
<name>OUT_3</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-63,169,-56.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>168.5,-63,169,-63</points>
<connection>
<GID>210</GID>
<name>ENABLE_0</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>153,-53.5,157.5,-53.5</points>
<connection>
<GID>209</GID>
<name>load</name></connection>
<intersection>153 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>153,-53.5,153,-51.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-53.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107.5,36,117.5,36</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<connection>
<GID>231</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>123.5,37,137.5,37</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-60.5,137,-59</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-59,137,-59</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-60.5,138,-58</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-58,138,-58</points>
<connection>
<GID>216</GID>
<name>OUT_1</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-60.5,139,-57</points>
<connection>
<GID>217</GID>
<name>IN_2</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-57,139,-57</points>
<connection>
<GID>216</GID>
<name>OUT_2</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-60.5,140,-56</points>
<connection>
<GID>217</GID>
<name>IN_3</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-56,140,-56</points>
<connection>
<GID>216</GID>
<name>OUT_3</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-62.5,142,-56</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>141.5,-62.5,142,-62.5</points>
<connection>
<GID>217</GID>
<name>ENABLE_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-53,130.5,-51</points>
<connection>
<GID>216</GID>
<name>load</name></connection>
<connection>
<GID>220</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-60.5,110,-59</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-59,110,-59</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-60.5,111,-58</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-58,111,-58</points>
<connection>
<GID>223</GID>
<name>OUT_1</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-60.5,112,-57</points>
<connection>
<GID>224</GID>
<name>IN_2</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-57,112,-57</points>
<connection>
<GID>223</GID>
<name>OUT_2</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-60.5,113,-56</points>
<connection>
<GID>224</GID>
<name>IN_3</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-56,113,-56</points>
<connection>
<GID>223</GID>
<name>OUT_3</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-62.5,115,-56</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-62.5,115,-62.5</points>
<connection>
<GID>224</GID>
<name>ENABLE_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>103.5,-53,103.5,-51</points>
<connection>
<GID>223</GID>
<name>load</name></connection>
<connection>
<GID>227</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,103.5,116.5,103.5</points>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<connection>
<GID>249</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>122.5,104.5,136.5,104.5</points>
<connection>
<GID>247</GID>
<name>OUT</name></connection>
<connection>
<GID>250</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>123.5,74,137,74</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<connection>
<GID>254</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,38,112,77</points>
<intersection>38 22</intersection>
<intersection>45.5 9</intersection>
<intersection>52 10</intersection>
<intersection>59 6</intersection>
<intersection>67.5 4</intersection>
<intersection>75 1</intersection>
<intersection>77 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,75,117.5,75</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106.5,77,112,77</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>112,67.5,117.5,67.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>112,59,117.5,59</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>112,45.5,117.5,45.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>112,52,117.5,52</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>112,38,117.5,38</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,72,115,73</points>
<intersection>72 2</intersection>
<intersection>73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,73,117.5,73</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107,72,115,72</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107.5,65.5,117.5,65.5</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<connection>
<GID>257</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>123.5,66.5,137.5,66.5</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<connection>
<GID>258</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194,99,229.5,99</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>261</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>51,-2.5,61.5,-2.5</points>
<connection>
<GID>50</GID>
<name>IN_3</name></connection>
<intersection>51 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>51,-2.5,51,-1</points>
<connection>
<GID>24</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-2.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,11.5,43,18</points>
<connection>
<GID>54</GID>
<name>count_enable</name></connection>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,14.5,2.5,15.5</points>
<intersection>14.5 2</intersection>
<intersection>15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,15.5,7,15.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,14.5,2.5,14.5</points>
<connection>
<GID>49</GID>
<name>OUT_2</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,12.5,3.5,13.5</points>
<intersection>12.5 1</intersection>
<intersection>13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,12.5,7,12.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,13.5,3.5,13.5</points>
<connection>
<GID>49</GID>
<name>OUT_1</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,0.5,112,18</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,0.5,112,0.5</points>
<connection>
<GID>62</GID>
<name>OUT_6</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,1.5,110,18.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>1.5 1</intersection>
<intersection>11 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,1.5,110,1.5</points>
<connection>
<GID>62</GID>
<name>OUT_7</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>110,11,133.5,11</points>
<connection>
<GID>360</GID>
<name>ENABLE</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,11.5,42,19.5</points>
<connection>
<GID>54</GID>
<name>load</name></connection>
<connection>
<GID>260</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-10.5,19.5,-10.5</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>15.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>15.5,-11,15.5,-10.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-7,21.5,-5</points>
<connection>
<GID>305</GID>
<name>SEL_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-5,21.5,-5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-8.5,19.5,-8.5</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<connection>
<GID>307</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-10,25,-9.5</points>
<intersection>-10 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-10,27.5,-10</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-9.5,25,-9.5</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-16,25.5,-12</points>
<connection>
<GID>309</GID>
<name>OUT</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-12,27.5,-12</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-15,15.5,-14</points>
<intersection>-15 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-15,19.5,-15</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-14,15.5,-14</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-17.5,16,-17</points>
<intersection>-17.5 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-17,19.5,-17</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-17.5,16,-17.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-11,42,0.5</points>
<connection>
<GID>54</GID>
<name>clock</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-11,42,-11</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-13.5,-8.5,-11.5,-8.5</points>
<connection>
<GID>317</GID>
<name>Q</name></connection>
<connection>
<GID>315</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20.5,-10.5,-19.5,-10.5</points>
<connection>
<GID>317</GID>
<name>clock</name></connection>
<intersection>-20.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-20.5,-14,-20.5,-10.5</points>
<intersection>-14 10</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-33.5,-14,-20.5,-14</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>-20.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>12</ID>
<points>-21.5,-12.5,-19.5,-12.5</points>
<connection>
<GID>317</GID>
<name>K</name></connection>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,-8.5,-19.5,-8.5</points>
<connection>
<GID>317</GID>
<name>J</name></connection>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<intersection>-26 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-26,-12.5,-26,-8.5</points>
<intersection>-12.5 17</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-26,-12.5,-25.5,-12.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>-26 14</intersection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-65,55.5,-65</points>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<intersection>34.5 16</intersection>
<intersection>35.5 17</intersection>
<intersection>36.5 18</intersection>
<intersection>43 19</intersection>
<intersection>44 20</intersection>
<intersection>45 10</intersection>
<intersection>51.5 5</intersection>
<intersection>52.5 6</intersection>
<intersection>53.5 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>51.5,-67,51.5,-65</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>-65 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>52.5,-67,52.5,-65</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<intersection>-65 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>53.5,-67,53.5,-65</points>
<connection>
<GID>349</GID>
<name>IN_2</name></connection>
<intersection>-65 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>45,-67,45,-65</points>
<connection>
<GID>348</GID>
<name>IN_2</name></connection>
<intersection>-65 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>34.5,-67,34.5,-65</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>-65 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>35.5,-67,35.5,-65</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>-65 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>36.5,-67,36.5,-65</points>
<connection>
<GID>347</GID>
<name>IN_2</name></connection>
<intersection>-65 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>43,-67,43,-65</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>-65 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>44,-67,44,-65</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<intersection>-65 1</intersection></vsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-64,40.5,-62</points>
<connection>
<GID>327</GID>
<name>A_less_B</name></connection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-64,54.5,-64</points>
<intersection>40.5 0</intersection>
<intersection>54.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-67,54.5,-64</points>
<connection>
<GID>349</GID>
<name>IN_3</name></connection>
<intersection>-64 2</intersection></vsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-66,39.5,-60</points>
<intersection>-66 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-60,40.5,-60</points>
<connection>
<GID>327</GID>
<name>A_equal_B</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-66,46,-66</points>
<intersection>39.5 0</intersection>
<intersection>46 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46,-67,46,-66</points>
<connection>
<GID>348</GID>
<name>IN_3</name></connection>
<intersection>-66 2</intersection></vsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-67,37.5,-58</points>
<connection>
<GID>347</GID>
<name>IN_3</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-58,40.5,-58</points>
<connection>
<GID>327</GID>
<name>A_greater_B</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-86,40,-69</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-69,40,-69</points>
<connection>
<GID>347</GID>
<name>ENABLE_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-86,48.5,-69</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-69,48.5,-69</points>
<connection>
<GID>348</GID>
<name>ENABLE_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-86,58,-69</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-69,58,-69</points>
<connection>
<GID>349</GID>
<name>ENABLE_0</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177.5,100,177.5,103.5</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177.5,100,188,100</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>177.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,49.5,158.5,104.5</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>49.5 3</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158.5,58,175.5,58</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>158.5,49.5,230,49.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,42,155.5,104.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>42 5</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,56,175.5,56</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>155.5,42,230,42</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,46,153,104.5</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>46 5</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153,54,175.5,54</points>
<connection>
<GID>380</GID>
<name>IN_2</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>153,46,230,46</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>181.5,56,197.5,56</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<intersection>197.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>197.5,56,197.5,85.5</points>
<intersection>56 1</intersection>
<intersection>85.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>197.5,85.5,198.5,85.5</points>
<connection>
<GID>395</GID>
<name>IN_1</name></connection>
<intersection>197.5 3</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-42.9134,2207.06,1735.09,1298.06</PageViewport></page 1>
<page 2>
<PageViewport>-42.9134,2207.06,1735.09,1298.06</PageViewport></page 2>
<page 3>
<PageViewport>-42.9134,2207.06,1735.09,1298.06</PageViewport></page 3>
<page 4>
<PageViewport>-42.9134,2207.06,1735.09,1298.06</PageViewport></page 4>
<page 5>
<PageViewport>-42.9134,2207.06,1735.09,1298.06</PageViewport></page 5>
<page 6>
<PageViewport>-42.9134,2207.06,1735.09,1298.06</PageViewport></page 6>
<page 7>
<PageViewport>-42.9134,2207.06,1735.09,1298.06</PageViewport></page 7>
<page 8>
<PageViewport>-42.9134,2207.06,1735.09,1298.06</PageViewport></page 8>
<page 9>
<PageViewport>-42.9134,2207.06,1735.09,1298.06</PageViewport></page 9></circuit>